TopicCode|ShortDesc|Desc
ENG01|Professional Sports on TV.|Do either of you have a favorite TV sport? How many hours per week do you spend watching it and other sporting events on TV?
ENG02|Pets.|Do either of you have a pet? If so, how much time each day do you spend with your pet? How important is your pet to you? 
ENG03|Life Partners.|What do each of you think is the most important thing to look for in a life partner? 
ENG04|Minimum Wage.|Do each of you feel the minimum wage increase - to <<$5.15 an hour - is sufficient? 
ENG05|Comedy.|How do you each draw the line between acceptable humor and humor that is in bad taste? 
ENG06|Hypothetical Situations. Perjury.|Do either of you think that you would commit perjury for a close friend or family member? 
ENG07|Hypothetical Situations. One Million Dollars to leave the US.|Would either of you accept one million dollars to leave the US and never return? If you were willing to leave, where would you go, what would you do? What would you miss the most about the US? What would you not miss? 
ENG08|Hypothetical Situations. Opening your own business|If each of you could open your own business, and money were not an issue, what type of business would you open? How would you go about doing this? Do you feel you would be a successful business owner? 
ENG09|Hypothetical Situations. Time Travel.|If each of you had the opportunity to go back in time and change something that you had done, what would it be and why? 
ENG10|Hypothetical Situations. An Anonymous Benefactor|If an unknown benefactor offered each of you a million dollars - with the only stipulation being that you could never speak to your best friend again - would you take the million dollars? 
ENG11|US Public Schools.|In your opinions, is there currently something seriously wrong with the public school system in the US, and if so, what can be done to correct it? 
ENG12|Affirmative Action.|Do either of you think affirmative action in hiring and promotion within the business community is a good policy? 
ENG13|Movies.|Do each of you enjoy going to the movies in a theater, or would you rather rent a movie and stay home? What was the last movie that you saw? Was it good or bad and why? 
ENG14|Computer games.|Do either of you play computer games? Do you play these games on the internet or on CD- ROM? What is your favorite game? 
ENG15|Current Events.|How do both of you keep up with current events? Do you get most of your news from TV, radio, newspapers, or people you know? 
ENG16|Hobbies.|What are your favorite hobbies? How much time do each of you spend pursuing your hobbies? Do you feel that every person needs at least one hobby? 
ENG17|Smoking. |How do you both feel about the movement to ban smoking in all public places? Do either of you think Smoking Prevention Programs, Counter-smoking ads, Help Quit hotlines and so on, are a good idea? 
ENG18|Terrorism.|Do you think most people would remain calm, or panic during a terrorist attack? How do you think each of you would react? 
ENG19|Televised Criminal Trials.|Do either of you feel that criminal trials, especially those involving high-profile individuals, should be televised? Have you ever watched any high-profile trials on TV? 
ENG20|Drug testing.|How do each of you feel about the practice of companies testing employees for drugs? Do you feel unannounced spot-checking for drugs to be an invasion of a person's privacy? 
ENG21|Family Values.|Do either of you feel that the increase in the divorce rate in the US has altered your behavior? Has it changed your views on the institution of marriage? 
ENG22|Censorship.|Do either of you think public or private schools have the right to forbid students to read certain books? 
ENG23|Health and Fitness.|Do each of you exercise regularly to maintain your health or fitness level? If so, what do you do? If not, would you like to start? 
ENG24|September 11.|What changes, if any, have either of you made in your life since the terrorist attacks of Sept 11, 2001? 
ENG25|Strikes by Professional Athletes.|How do each of you feel about the recent strikes by professional athletes? Do you think that professional athletes deserve the high salaries they currently receive? 
ENG26|Airport Security.|Do either of you think that heightened airport security lessens the chance of terrorist incidents in the air? 
ENG27|Issues in the Middle East. |What does each of you think about the current unrest in the Middle East? Do you feel that peace will ever be attained in the area? Should the US remain involved in the peace process? 
ENG28|Foreign Relations.|Do either of you consider any other countries to be a threat to US safety? If so, which countries and why? 
ENG29|Education.|What do each of you think about computers in education? Do they improve or harm education? 
ENG30|Family.|What does the word family mean to each of you? 
ENG31|Corporate Conduct in the US.|What do each of you think the government can do to curb illegal business activity? Has the cascade of corporate scandals caused the mild recession and decline in the US stock market and economy? How have the scandals affected you? 
ENG32|Outdoor Activities.|Do you like cold weather or warm weather activities the best? Do you like outside or inside activities better? Each of you should talk about your favorite activities. 
ENG33|Friends.|Are either of you the type of person who has lots of friends and acquaintances or do you just have a few close friends? Each of you should talk about your best friend or friends. 
ENG34|Food.|Which do each of you like better--eating at a restaurant or at home? Describe your perfect meal. 
ENG35|Illness.|When the seasons change, many people get ill. Do either of you? What do you do to keep yourself well? There is a saying, "A cold lasts seven days if you don't go to the doctor and a week if you do." Do you both agree? 
ENG36|Personal Habits.|According to each of you, which is worse: gossiping, smoking, drinking alcohol or caffeine excessively, overeating, or not exercising? 
ENG37|Reality TV.|Do either of you watch reality shows on TV. If so, which one or ones? Why do you think that reality based television programming, shows like "Survivor" or "Who Wants to Marry a Millionaire" are so popular? 
ENG38|Arms Inspections in Iraq.|What, if anything, do you both think the US should do about Iraq? Do you think that disarming Iraq should be a major priority for the US? 
ENG39|Holidays.|Do either of you have a favorit holiday? Why? If either of you you could create a holiday, what would it be and how would you have people celebrate it? 
ENG40|Bioterrorism.|What do you both think the US can do to prevent a bioterrorist attack? 
